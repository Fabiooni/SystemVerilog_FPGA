--------------------------------------------------------------------------------
--                     FixRealKCM_comb_uid6_T0_comb_uid9
-- VHDL generated for Virtex6 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: 0.000000ns
--  approx. output signal timings: Y: 0.655000ns

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_comb_uid6_T0_comb_uid9 is
    port (X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(9 downto 0)   );
end entity;

architecture arch of FixRealKCM_comb_uid6_T0_comb_uid9 is
signal Y0 :  std_logic_vector(9 downto 0);
   -- timing of Y0: 0.655000ns
signal Y1 :  std_logic_vector(9 downto 0);
   -- timing of Y1: 0.655000ns
begin
   with X  select  Y0 <= 
      "0000000000" when "000000",
      "0000001101" when "000001",
      "0000011001" when "000010",
      "0000100110" when "000011",
      "0000110010" when "000100",
      "0000111111" when "000101",
      "0001001011" when "000110",
      "0001011000" when "000111",
      "0001100101" when "001000",
      "0001110001" when "001001",
      "0001111110" when "001010",
      "0010001010" when "001011",
      "0010010111" when "001100",
      "0010100011" when "001101",
      "0010110000" when "001110",
      "0010111100" when "001111",
      "0011001001" when "010000",
      "0011010110" when "010001",
      "0011100010" when "010010",
      "0011101111" when "010011",
      "0011111011" when "010100",
      "0100001000" when "010101",
      "0100010100" when "010110",
      "0100100001" when "010111",
      "0100101110" when "011000",
      "0100111010" when "011001",
      "0101000111" when "011010",
      "0101010011" when "011011",
      "0101100000" when "011100",
      "0101101100" when "011101",
      "0101111001" when "011110",
      "0110000110" when "011111",
      "0110010010" when "100000",
      "0110011111" when "100001",
      "0110101011" when "100010",
      "0110111000" when "100011",
      "0111000100" when "100100",
      "0111010001" when "100101",
      "0111011110" when "100110",
      "0111101010" when "100111",
      "0111110111" when "101000",
      "1000000011" when "101001",
      "1000010000" when "101010",
      "1000011100" when "101011",
      "1000101001" when "101100",
      "1000110101" when "101101",
      "1001000010" when "101110",
      "1001001111" when "101111",
      "1001011011" when "110000",
      "1001101000" when "110001",
      "1001110100" when "110010",
      "1010000001" when "110011",
      "1010001101" when "110100",
      "1010011010" when "110101",
      "1010100111" when "110110",
      "1010110011" when "110111",
      "1011000000" when "111000",
      "1011001100" when "111001",
      "1011011001" when "111010",
      "1011100101" when "111011",
      "1011110010" when "111100",
      "1011111111" when "111101",
      "1100001011" when "111110",
      "1100011000" when "111111",
      "----------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                     FixRealKCM_comb_uid6_T1_comb_uid11
-- VHDL generated for Virtex6 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: 0.000000ns
--  approx. output signal timings: Y: 0.649000ns

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_comb_uid6_T1_comb_uid11 is
    port (X : in  std_logic_vector(1 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of FixRealKCM_comb_uid6_T1_comb_uid11 is
signal Y0 :  std_logic_vector(3 downto 0);
   -- timing of Y0: 0.649000ns
signal Y1 :  std_logic_vector(3 downto 0);
   -- timing of Y1: 0.649000ns
begin
   with X  select  Y0 <= 
      "0000" when "00",
      "0011" when "01",
      "0110" when "10",
      "1001" when "11",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           SinCosTable_comb_uid4
-- VHDL generated for Virtex6 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: 0.366000ns
--  approx. output signal timings: Y: 2.236000ns

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity SinCosTable_comb_uid4 is
    port (X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(39 downto 0)   );
end entity;

architecture arch of SinCosTable_comb_uid4 is
signal Y0 :  std_logic_vector(39 downto 0);
   -- timing of Y0: 2.236000ns
signal Y1 :  std_logic_vector(39 downto 0);
   -- timing of Y1: 2.236000ns
begin
   with X  select  Y0 <= 
      "0000000000000000100011111111111111111000" when "0000000000",
      "0000000000110010110011111111111111111000" when "0000000001",
      "0000000001100101000011111111111111110111" when "0000000010",
      "0000000010010111010111111111111111110101" when "0000000011",
      "0000000011001001100111111111111111110011" when "0000000100",
      "0000000011111011110111111111111111110000" when "0000000101",
      "0000000100101110000111111111111111101101" when "0000000110",
      "0000000101100000011011111111111111101001" when "0000000111",
      "0000000110010010101011111111111111100100" when "0000001000",
      "0000000111000100111011111111111111011111" when "0000001001",
      "0000000111110111001011111111111111011001" when "0000001010",
      "0000001000101001011011111111111111010011" when "0000001011",
      "0000001001011011101111111111111111001100" when "0000001100",
      "0000001010001101111111111111111111000100" when "0000001101",
      "0000001011000000001111111111111110111100" when "0000001110",
      "0000001011110010011111111111111110110011" when "0000001111",
      "0000001100100100101111111111111110101001" when "0000010000",
      "0000001101010111000011111111111110011111" when "0000010001",
      "0000001110001001010011111111111110010100" when "0000010010",
      "0000001110111011100011111111111110001001" when "0000010011",
      "0000001111101101110011111111111101111101" when "0000010100",
      "0000010000100000000011111111111101110000" when "0000010101",
      "0000010001010010010011111111111101100011" when "0000010110",
      "0000010010000100100011111111111101010101" when "0000010111",
      "0000010010110110110111111111111101000110" when "0000011000",
      "0000010011101001000111111111111100110111" when "0000011001",
      "0000010100011011010111111111111100101000" when "0000011010",
      "0000010101001101100111111111111100010111" when "0000011011",
      "0000010101111111110111111111111100000110" when "0000011100",
      "0000010110110010000111111111111011110101" when "0000011101",
      "0000010111100100010111111111111011100010" when "0000011110",
      "0000011000010110100111111111111011010000" when "0000011111",
      "0000011001001000110111111111111010111100" when "0000100000",
      "0000011001111011000111111111111010101000" when "0000100001",
      "0000011010101101010111111111111010010011" when "0000100010",
      "0000011011011111100111111111111001111110" when "0000100011",
      "0000011100010001110111111111111001101000" when "0000100100",
      "0000011101000100000111111111111001010010" when "0000100101",
      "0000011101110110010111111111111000111011" when "0000100110",
      "0000011110101000100111111111111000100011" when "0000100111",
      "0000011111011010110011111111111000001011" when "0000101000",
      "0000100000001101000011111111110111110010" when "0000101001",
      "0000100000111111010011111111110111011000" when "0000101010",
      "0000100001110001100011111111110110111110" when "0000101011",
      "0000100010100011110011111111110110100011" when "0000101100",
      "0000100011010101111111111111110110001000" when "0000101101",
      "0000100100001000001111111111110101101011" when "0000101110",
      "0000100100111010011111111111110101001111" when "0000101111",
      "0000100101101100101111111111110100110001" when "0000110000",
      "0000100110011110111011111111110100010100" when "0000110001",
      "0000100111010001001011111111110011110101" when "0000110010",
      "0000101000000011011011111111110011010110" when "0000110011",
      "0000101000110101100111111111110010110110" when "0000110100",
      "0000101001100111110111111111110010010110" when "0000110101",
      "0000101010011010000011111111110001110101" when "0000110110",
      "0000101011001100010011111111110001010011" when "0000110111",
      "0000101011111110011111111111110000110001" when "0000111000",
      "0000101100110000101111111111110000001110" when "0000111001",
      "0000101101100010111011111111101111101011" when "0000111010",
      "0000101110010101001011111111101111000111" when "0000111011",
      "0000101111000111010111111111101110100010" when "0000111100",
      "0000101111111001100011111111101101111101" when "0000111101",
      "0000110000101011110011111111101101010111" when "0000111110",
      "0000110001011101111111111111101100110000" when "0000111111",
      "0000110010010000001011111111101100001001" when "0001000000",
      "0000110011000010011011111111101011100001" when "0001000001",
      "0000110011110100100111111111101010111001" when "0001000010",
      "0000110100100110110011111111101010010000" when "0001000011",
      "0000110101011000111111111111101001100110" when "0001000100",
      "0000110110001011001011111111101000111100" when "0001000101",
      "0000110110111101010111111111101000010001" when "0001000110",
      "0000110111101111100011111111100111100110" when "0001000111",
      "0000111000100001110011111111100110111010" when "0001001000",
      "0000111001010011111111111111100110001101" when "0001001001",
      "0000111010000110000111111111100101100000" when "0001001010",
      "0000111010111000010011111111100100110010" when "0001001011",
      "0000111011101010011111111111100100000011" when "0001001100",
      "0000111100011100101011111111100011010100" when "0001001101",
      "0000111101001110110111111111100010100100" when "0001001110",
      "0000111110000001000011111111100001110100" when "0001001111",
      "0000111110110011001011111111100001000011" when "0001010000",
      "0000111111100101010111111111100000010001" when "0001010001",
      "0001000000010111100011111111011111011111" when "0001010010",
      "0001000001001001101011111111011110101100" when "0001010011",
      "0001000001111011110111111111011101111001" when "0001010100",
      "0001000010101110000011111111011101000100" when "0001010101",
      "0001000011100000001011111111011100010000" when "0001010110",
      "0001000100010010010111111111011011011010" when "0001010111",
      "0001000101000100011111111111011010100100" when "0001011000",
      "0001000101110110100111111111011001101110" when "0001011001",
      "0001000110101000110011111111011000110111" when "0001011010",
      "0001000111011010111011111111010111111111" when "0001011011",
      "0001001000001101000011111111010111000111" when "0001011100",
      "0001001000111111001011111111010110001110" when "0001011101",
      "0001001001110001010111111111010101010100" when "0001011110",
      "0001001010100011011111111111010100011010" when "0001011111",
      "0001001011010101100111111111010011011111" when "0001100000",
      "0001001100000111101111111111010010100011" when "0001100001",
      "0001001100111001110111111111010001100111" when "0001100010",
      "0001001101101011111111111111010000101011" when "0001100011",
      "0001001110011110000111111111001111101101" when "0001100100",
      "0001001111010000001111111111001110101111" when "0001100101",
      "0001010000000010010011111111001101110001" when "0001100110",
      "0001010000110100011011111111001100110010" when "0001100111",
      "0001010001100110100011111111001011110010" when "0001101000",
      "0001010010011000100111111111001010110010" when "0001101001",
      "0001010011001010101111111111001001110000" when "0001101010",
      "0001010011111100110111111111001000101111" when "0001101011",
      "0001010100101110111011111111000111101101" when "0001101100",
      "0001010101100001000011111111000110101010" when "0001101101",
      "0001010110010011000111111111000101100110" when "0001101110",
      "0001010111000101001011111111000100100010" when "0001101111",
      "0001010111110111010011111111000011011110" when "0001110000",
      "0001011000101001010111111111000010011000" when "0001110001",
      "0001011001011011011011111111000001010010" when "0001110010",
      "0001011010001101011111111111000000001100" when "0001110011",
      "0001011010111111100011111110111111000101" when "0001110100",
      "0001011011110001100111111110111101111101" when "0001110101",
      "0001011100100011101011111110111100110100" when "0001110110",
      "0001011101010101101111111110111011101011" when "0001110111",
      "0001011110000111110011111110111010100010" when "0001111000",
      "0001011110111001110111111110111001011000" when "0001111001",
      "0001011111101011111011111110111000001101" when "0001111010",
      "0001100000011101111011111110110111000001" when "0001111011",
      "0001100001001111111111111110110101110101" when "0001111100",
      "0001100010000001111111111110110100101001" when "0001111101",
      "0001100010110100000011111110110011011011" when "0001111110",
      "0001100011100110000011111110110010001101" when "0001111111",
      "0001100100011000000111111110110000111111" when "0010000000",
      "0001100101001010000111111110101111110000" when "0010000001",
      "0001100101111100000111111110101110100000" when "0010000010",
      "0001100110101110001011111110101101010000" when "0010000011",
      "0001100111100000001011111110101011111111" when "0010000100",
      "0001101000010010001011111110101010101101" when "0010000101",
      "0001101001000100001011111110101001011011" when "0010000110",
      "0001101001110110001011111110101000001000" when "0010000111",
      "0001101010101000001011111110100110110101" when "0010001000",
      "0001101011011010001011111110100101100001" when "0010001001",
      "0001101100001100000111111110100100001100" when "0010001010",
      "0001101100111110000111111110100010110111" when "0010001011",
      "0001101101110000000111111110100001100001" when "0010001100",
      "0001101110100010000011111110100000001010" when "0010001101",
      "0001101111010100000011111110011110110011" when "0010001110",
      "0001110000000101111111111110011101011011" when "0010001111",
      "0001110000110111111111111110011100000011" when "0010010000",
      "0001110001101001111011111110011010101010" when "0010010001",
      "0001110010011011110111111110011001010001" when "0010010010",
      "0001110011001101110011111110010111110110" when "0010010011",
      "0001110011111111101111111110010110011100" when "0010010100",
      "0001110100110001101011111110010101000000" when "0010010101",
      "0001110101100011100111111110010011100100" when "0010010110",
      "0001110110010101100011111110010010001000" when "0010010111",
      "0001110111000111011111111110010000101010" when "0010011000",
      "0001110111111001011011111110001111001100" when "0010011001",
      "0001111000101011010011111110001101101110" when "0010011010",
      "0001111001011101001111111110001100001111" when "0010011011",
      "0001111010001111001011111110001010101111" when "0010011100",
      "0001111011000001000011111110001001001111" when "0010011101",
      "0001111011110010111011111110000111101110" when "0010011110",
      "0001111100100100110111111110000110001100" when "0010011111",
      "0001111101010110101111111110000100101010" when "0010100000",
      "0001111110001000100111111110000011001000" when "0010100001",
      "0001111110111010011111111110000001100100" when "0010100010",
      "0001111111101100010111111110000000000000" when "0010100011",
      "0010000000011110001111111101111110011100" when "0010100100",
      "0010000001010000000111111101111100110110" when "0010100101",
      "0010000010000001111111111101111011010001" when "0010100110",
      "0010000010110011110011111101111001101010" when "0010100111",
      "0010000011100101101011111101111000000011" when "0010101000",
      "0010000100010111100011111101110110011100" when "0010101001",
      "0010000101001001010111111101110100110011" when "0010101010",
      "0010000101111011001011111101110011001010" when "0010101011",
      "0010000110101101000011111101110001100001" when "0010101100",
      "0010000111011110110111111101101111110111" when "0010101101",
      "0010001000010000101011111101101110001100" when "0010101110",
      "0010001001000010011111111101101100100001" when "0010101111",
      "0010001001110100010011111101101010110101" when "0010110000",
      "0010001010100110000111111101101001001000" when "0010110001",
      "0010001011010111111011111101100111011011" when "0010110010",
      "0010001100001001101011111101100101101101" when "0010110011",
      "0010001100111011011111111101100011111111" when "0010110100",
      "0010001101101101001111111101100010010000" when "0010110101",
      "0010001110011111000011111101100000100000" when "0010110110",
      "0010001111010000110011111101011110110000" when "0010110111",
      "0010010000000010100111111101011100111111" when "0010111000",
      "0010010000110100010111111101011011001110" when "0010111001",
      "0010010001100110000111111101011001011100" when "0010111010",
      "0010010010010111110111111101010111101001" when "0010111011",
      "0010010011001001100111111101010101110110" when "0010111100",
      "0010010011111011010111111101010100000010" when "0010111101",
      "0010010100101101000011111101010010001110" when "0010111110",
      "0010010101011110110011111101010000011001" when "0010111111",
      "0010010110010000100011111101001110100011" when "0011000000",
      "0010010111000010001111111101001100101101" when "0011000001",
      "0010010111110011111111111101001010110110" when "0011000010",
      "0010011000100101101011111101001000111110" when "0011000011",
      "0010011001010111010111111101000111000110" when "0011000100",
      "0010011010001001000011111101000101001101" when "0011000101",
      "0010011010111010101111111101000011010100" when "0011000110",
      "0010011011101100011011111101000001011010" when "0011000111",
      "0010011100011110000111111100111111011111" when "0011001000",
      "0010011101001111110011111100111101100100" when "0011001001",
      "0010011110000001011011111100111011101000" when "0011001010",
      "0010011110110011000111111100111001101100" when "0011001011",
      "0010011111100100101111111100110111101111" when "0011001100",
      "0010100000010110011011111100110101110001" when "0011001101",
      "0010100001001000000011111100110011110011" when "0011001110",
      "0010100001111001101011111100110001110100" when "0011001111",
      "0010100010101011010011111100101111110101" when "0011010000",
      "0010100011011100111011111100101101110101" when "0011010001",
      "0010100100001110100011111100101011110100" when "0011010010",
      "0010100101000000001011111100101001110011" when "0011010011",
      "0010100101110001110011111100100111110001" when "0011010100",
      "0010100110100011010111111100100101101110" when "0011010101",
      "0010100111010100111111111100100011101011" when "0011010110",
      "0010101000000110100011111100100001101000" when "0011010111",
      "0010101000111000000111111100011111100011" when "0011011000",
      "0010101001101001101011111100011101011110" when "0011011001",
      "0010101010011011010011111100011011011001" when "0011011010",
      "0010101011001100110111111100011001010011" when "0011011011",
      "0010101011111110010111111100010111001100" when "0011011100",
      "0010101100101111111011111100010101000100" when "0011011101",
      "0010101101100001011111111100010010111100" when "0011011110",
      "0010101110010010111111111100010000110100" when "0011011111",
      "0010101111000100100011111100001110101011" when "0011100000",
      "0010101111110110000011111100001100100001" when "0011100001",
      "0010110000100111100011111100001010010111" when "0011100010",
      "0010110001011001000111111100001000001100" when "0011100011",
      "0010110010001010100111111100000110000000" when "0011100100",
      "0010110010111100000011111100000011110100" when "0011100101",
      "0010110011101101100011111100000001100111" when "0011100110",
      "0010110100011111000011111011111111011001" when "0011100111",
      "0010110101010000100011111011111101001011" when "0011101000",
      "0010110110000001111111111011111010111101" when "0011101001",
      "0010110110110011011011111011111000101101" when "0011101010",
      "0010110111100100111011111011110110011110" when "0011101011",
      "0010111000010110010111111011110100001101" when "0011101100",
      "0010111001000111110011111011110001111100" when "0011101101",
      "0010111001111001001111111011101111101010" when "0011101110",
      "0010111010101010101011111011101101011000" when "0011101111",
      "0010111011011100000011111011101011000101" when "0011110000",
      "0010111100001101011111111011101000110010" when "0011110001",
      "0010111100111110110111111011100110011101" when "0011110010",
      "0010111101110000010011111011100100001001" when "0011110011",
      "0010111110100001101011111011100001110011" when "0011110100",
      "0010111111010011000011111011011111011101" when "0011110101",
      "0011000000000100011011111011011101000111" when "0011110110",
      "0011000000110101110011111011011010110000" when "0011110111",
      "0011000001100111001011111011011000011000" when "0011111000",
      "0011000010011000100011111011010110000000" when "0011111001",
      "0011000011001001110111111011010011100111" when "0011111010",
      "0011000011111011001111111011010001001101" when "0011111011",
      "0011000100101100100011111011001110110011" when "0011111100",
      "0011000101011101110111111011001100011000" when "0011111101",
      "0011000110001111001011111011001001111101" when "0011111110",
      "0011000111000000011111111011000111100001" when "0011111111",
      "0011000111110001110011111011000101000100" when "0100000000",
      "0011001000100011000111111011000010100111" when "0100000001",
      "0011001001010100010111111011000000001001" when "0100000010",
      "0011001010000101101011111010111101101011" when "0100000011",
      "0011001010110110111011111010111011001100" when "0100000100",
      "0011001011101000001011111010111000101100" when "0100000101",
      "0011001100011001011011111010110110001100" when "0100000110",
      "0011001101001010101011111010110011101011" when "0100000111",
      "0011001101111011111011111010110001001010" when "0100001000",
      "0011001110101101001011111010101110101000" when "0100001001",
      "0011001111011110011011111010101100000101" when "0100001010",
      "0011010000001111100111111010101001100010" when "0100001011",
      "0011010001000000110011111010100110111110" when "0100001100",
      "0011010001110010000011111010100100011001" when "0100001101",
      "0011010010100011001111111010100001110100" when "0100001110",
      "0011010011010100011011111010011111001111" when "0100001111",
      "0011010100000101100111111010011100101000" when "0100010000",
      "0011010100110110101111111010011010000010" when "0100010001",
      "0011010101100111111011111010010111011010" when "0100010010",
      "0011010110011001000111111010010100110010" when "0100010011",
      "0011010111001010001111111010010010001001" when "0100010100",
      "0011010111111011010111111010001111100000" when "0100010101",
      "0011011000101100011111111010001100110110" when "0100010110",
      "0011011001011101100111111010001010001100" when "0100010111",
      "0011011010001110101111111010000111100001" when "0100011000",
      "0011011010111111110111111010000100110101" when "0100011001",
      "0011011011110000111011111010000010001001" when "0100011010",
      "0011011100100010000011111001111111011100" when "0100011011",
      "0011011101010011000111111001111100101110" when "0100011100",
      "0011011110000100001011111001111010000000" when "0100011101",
      "0011011110110101001111111001110111010001" when "0100011110",
      "0011011111100110010011111001110100100010" when "0100011111",
      "0011100000010111010111111001110001110010" when "0100100000",
      "0011100001001000010111111001101111000010" when "0100100001",
      "0011100001111001011011111001101100010001" when "0100100010",
      "0011100010101010011011111001101001011111" when "0100100011",
      "0011100011011011011011111001100110101101" when "0100100100",
      "0011100100001100011111111001100011111010" when "0100100101",
      "0011100100111101011111111001100001000110" when "0100100110",
      "0011100101101110011011111001011110010010" when "0100100111",
      "0011100110011111011011111001011011011101" when "0100101000",
      "0011100111010000011011111001011000101000" when "0100101001",
      "0011101000000001010111111001010101110010" when "0100101010",
      "0011101000110010010011111001010010111100" when "0100101011",
      "0011101001100011001111111001010000000100" when "0100101100",
      "0011101010010100001011111001001101001101" when "0100101101",
      "0011101011000101000111111001001010010100" when "0100101110",
      "0011101011110110000011111001000111011011" when "0100101111",
      "0011101100100110111011111001000100100010" when "0100110000",
      "0011101101010111110111111001000001101000" when "0100110001",
      "0011101110001000101111111000111110101101" when "0100110010",
      "0011101110111001100111111000111011110010" when "0100110011",
      "0011101111101010011111111000111000110110" when "0100110100",
      "0011110000011011010111111000110101111001" when "0100110101",
      "0011110001001100001111111000110010111100" when "0100110110",
      "0011110001111101000011111000101111111110" when "0100110111",
      "0011110010101101110111111000101101000000" when "0100111000",
      "0011110011011110101111111000101010000001" when "0100111001",
      "0011110100001111100011111000100111000010" when "0100111010",
      "0011110101000000010111111000100100000010" when "0100111011",
      "0011110101110001001011111000100001000001" when "0100111100",
      "0011110110100001111011111000011110000000" when "0100111101",
      "0011110111010010101111111000011010111110" when "0100111110",
      "0011111000000011011111111000010111111011" when "0100111111",
      "0011111000110100001111111000010100111000" when "0101000000",
      "0011111001100100111111111000010001110100" when "0101000001",
      "0011111010010101101111111000001110110000" when "0101000010",
      "0011111011000110011111111000001011101011" when "0101000011",
      "0011111011110111001111111000001000100110" when "0101000100",
      "0011111100100111111011111000000101011111" when "0101000101",
      "0011111101011000100111111000000010011001" when "0101000110",
      "0011111110001001010111110111111111010001" when "0101000111",
      "0011111110111010000011110111111100001010" when "0101001000",
      "0011111111101010101011110111111001000001" when "0101001001",
      "0100000000011011010111110111110101111000" when "0101001010",
      "0100000001001100000011110111110010101110" when "0101001011",
      "0100000001111100101011110111101111100100" when "0101001100",
      "0100000010101101010011110111101100011001" when "0101001101",
      "0100000011011101111011110111101001001110" when "0101001110",
      "0100000100001110100011110111100110000010" when "0101001111",
      "0100000100111111001011110111100010110101" when "0101010000",
      "0100000101101111110011110111011111101000" when "0101010001",
      "0100000110100000010111110111011100011010" when "0101010010",
      "0100000111010000111011110111011001001011" when "0101010011",
      "0100001000000001011111110111010101111100" when "0101010100",
      "0100001000110010000011110111010010101101" when "0101010101",
      "0100001001100010100111110111001111011100" when "0101010110",
      "0100001010010011001011110111001100001011" when "0101010111",
      "0100001011000011101011110111001000111010" when "0101011000",
      "0100001011110100001111110111000101101000" when "0101011001",
      "0100001100100100101111110111000010010101" when "0101011010",
      "0100001101010101001111110110111111000010" when "0101011011",
      "0100001110000101101111110110111011101110" when "0101011100",
      "0100001110110110001011110110111000011010" when "0101011101",
      "0100001111100110101011110110110101000101" when "0101011110",
      "0100010000010111000111110110110001101111" when "0101011111",
      "0100010001000111100011110110101110011001" when "0101100000",
      "0100010001110111111111110110101011000010" when "0101100001",
      "0100010010101000011011110110100111101011" when "0101100010",
      "0100010011011000110111110110100100010011" when "0101100011",
      "0100010100001001001111110110100000111010" when "0101100100",
      "0100010100111001101011110110011101100001" when "0101100101",
      "0100010101101010000011110110011010000111" when "0101100110",
      "0100010110011010011011110110010110101101" when "0101100111",
      "0100010111001010110011110110010011010010" when "0101101000",
      "0100010111111011001011110110001111110110" when "0101101001",
      "0100011000101011011111110110001100011010" when "0101101010",
      "0100011001011011110011110110001000111110" when "0101101011",
      "0100011010001100001011110110000101100000" when "0101101100",
      "0100011010111100011111110110000010000010" when "0101101101",
      "0100011011101100101111110101111110100100" when "0101101110",
      "0100011100011101000011110101111011000101" when "0101101111",
      "0100011101001101010111110101110111100101" when "0101110000",
      "0100011101111101100111110101110100000101" when "0101110001",
      "0100011110101101110111110101110000100100" when "0101110010",
      "0100011111011110000111110101101101000010" when "0101110011",
      "0100100000001110010111110101101001100000" when "0101110100",
      "0100100000111110100111110101100101111110" when "0101110101",
      "0100100001101110110011110101100010011010" when "0101110110",
      "0100100010011110111111110101011110110111" when "0101110111",
      "0100100011001111001011110101011011010010" when "0101111000",
      "0100100011111111010111110101010111101101" when "0101111001",
      "0100100100101111100011110101010100000111" when "0101111010",
      "0100100101011111101111110101010000100001" when "0101111011",
      "0100100110001111110111110101001100111010" when "0101111100",
      "0100100110111111111111110101001001010011" when "0101111101",
      "0100100111110000000111110101000101101011" when "0101111110",
      "0100101000100000001111110101000010000011" when "0101111111",
      "0100101001010000010111110100111110011001" when "0110000000",
      "0100101010000000011011110100111010110000" when "0110000001",
      "0100101010110000100011110100110111000101" when "0110000010",
      "0100101011100000100111110100110011011010" when "0110000011",
      "0100101100010000101011110100101111101111" when "0110000100",
      "0100101101000000101111110100101100000011" when "0110000101",
      "0100101101110000101111110100101000010110" when "0110000110",
      "0100101110100000110011110100100100101001" when "0110000111",
      "0100101111010000110011110100100000111011" when "0110001000",
      "0100110000000000110011110100011101001100" when "0110001001",
      "0100110000110000110011110100011001011101" when "0110001010",
      "0100110001100000110011110100010101101110" when "0110001011",
      "0100110010010000101111110100010001111101" when "0110001100",
      "0100110011000000101011110100001110001101" when "0110001101",
      "0100110011110000101011110100001010011011" when "0110001110",
      "0100110100100000100111110100000110101001" when "0110001111",
      "0100110101010000011111110100000010110111" when "0110010000",
      "0100110110000000011011110011111111000011" when "0110010001",
      "0100110110110000010011110011111011010000" when "0110010010",
      "0100110111100000001111110011110111011011" when "0110010011",
      "0100111000010000000111110011110011100110" when "0110010100",
      "0100111000111111111011110011101111110001" when "0110010101",
      "0100111001101111110011110011101011111011" when "0110010110",
      "0100111010011111101011110011101000000100" when "0110010111",
      "0100111011001111011111110011100100001101" when "0110011000",
      "0100111011111111010011110011100000010101" when "0110011001",
      "0100111100101111000111110011011100011100" when "0110011010",
      "0100111101011110110111110011011000100011" when "0110011011",
      "0100111110001110101011110011010100101010" when "0110011100",
      "0100111110111110011011110011010000101111" when "0110011101",
      "0100111111101110001011110011001100110101" when "0110011110",
      "0101000000011101111011110011001000111001" when "0110011111",
      "0101000001001101101011110011000100111101" when "0110100000",
      "0101000001111101011011110011000001000001" when "0110100001",
      "0101000010101101000111110010111101000100" when "0110100010",
      "0101000011011100110011110010111001000110" when "0110100011",
      "0101000100001100011111110010110101000111" when "0110100100",
      "0101000100111100001011110010110001001001" when "0110100101",
      "0101000101101011110011110010101101001001" when "0110100110",
      "0101000110011011011111110010101001001001" when "0110100111",
      "0101000111001011000111110010100101001000" when "0110101000",
      "0101000111111010101111110010100001000111" when "0110101001",
      "0101001000101010010111110010011101000101" when "0110101010",
      "0101001001011001111011110010011001000011" when "0110101011",
      "0101001010001001100011110010010101000000" when "0110101100",
      "0101001010111001000111110010010000111100" when "0110101101",
      "0101001011101000101011110010001100111000" when "0110101110",
      "0101001100011000001111110010001000110011" when "0110101111",
      "0101001101000111101111110010000100101110" when "0110110000",
      "0101001101110111010011110010000000101000" when "0110110001",
      "0101001110100110110011110001111100100010" when "0110110010",
      "0101001111010110010011110001111000011011" when "0110110011",
      "0101010000000101110011110001110100010011" when "0110110100",
      "0101010000110101001111110001110000001011" when "0110110101",
      "0101010001100100101111110001101100000010" when "0110110110",
      "0101010010010100001011110001100111111000" when "0110110111",
      "0101010011000011100111110001100011101110" when "0110111000",
      "0101010011110011000011110001011111100100" when "0110111001",
      "0101010100100010011011110001011011011001" when "0110111010",
      "0101010101010001110111110001010111001101" when "0110111011",
      "0101010110000001001111110001010011000001" when "0110111100",
      "0101010110110000100111110001001110110100" when "0110111101",
      "0101010111011111111011110001001010100110" when "0110111110",
      "0101011000001111010011110001000110011000" when "0110111111",
      "0101011000111110100111110001000010001001" when "0111000000",
      "0101011001101101111011110000111101111010" when "0111000001",
      "0101011010011101001111110000111001101010" when "0111000010",
      "0101011011001100100011110000110101011010" when "0111000011",
      "0101011011111011110011110000110001001001" when "0111000100",
      "0101011100101011000111110000101100110111" when "0111000101",
      "0101011101011010010111110000101000100101" when "0111000110",
      "0101011110001001100111110000100100010011" when "0111000111",
      "0101011110111000110011110000011111111111" when "0111001000",
      "0101011111101000000011110000011011101011" when "0111001001",
      "0101100000010111001111110000010111010111" when "0111001010",
      "0101100001000110011011110000010011000010" when "0111001011",
      "0101100001110101100111110000001110101100" when "0111001100",
      "0101100010100100101111110000001010010110" when "0111001101",
      "0101100011010011111011110000000101111111" when "0111001110",
      "0101100100000011000011110000000001101000" when "0111001111",
      "0101100100110010001011101111111101010000" when "0111010000",
      "0101100101100001010011101111111000111000" when "0111010001",
      "0101100110010000010111101111110100011111" when "0111010010",
      "0101100110111111011011101111110000000101" when "0111010011",
      "0101100111101110100011101111101011101011" when "0111010100",
      "0101101000011101100011101111100111010000" when "0111010101",
      "0101101001001100100111101111100010110101" when "0111010110",
      "0101101001111011100111101111011110011001" when "0111010111",
      "0101101010101010101011101111011001111100" when "0111011000",
      "0101101011011001101011101111010101011111" when "0111011001",
      "0101101100001000100111101111010001000001" when "0111011010",
      "0101101100110111100111101111001100100011" when "0111011011",
      "0101101101100110100011101111001000000100" when "0111011100",
      "0101101110010101100011101111000011100101" when "0111011101",
      "0101101111000100011011101110111111000101" when "0111011110",
      "0101101111110011010111101110111010100100" when "0111011111",
      "0101110000100010010011101110110110000011" when "0111100000",
      "0101110001010001001011101110110001100001" when "0111100001",
      "0101110010000000000011101110101100111111" when "0111100010",
      "0101110010101110111011101110101000011100" when "0111100011",
      "0101110011011101101111101110100011111001" when "0111100100",
      "0101110100001100100011101110011111010101" when "0111100101",
      "0101110100111011011011101110011010110000" when "0111100110",
      "0101110101101010001011101110010110001011" when "0111100111",
      "0101110110011000111111101110010001100101" when "0111101000",
      "0101110111000111110011101110001100111111" when "0111101001",
      "0101110111110110100011101110001000011000" when "0111101010",
      "0101111000100101010011101110000011110000" when "0111101011",
      "0101111001010100000011101101111111001000" when "0111101100",
      "0101111010000010101111101101111010100000" when "0111101101",
      "0101111010110001011011101101110101110110" when "0111101110",
      "0101111011100000001011101101110001001101" when "0111101111",
      "0101111100001110110011101101101100100010" when "0111110000",
      "0101111100111101011111101101100111110111" when "0111110001",
      "0101111101101100000111101101100011001100" when "0111110010",
      "0101111110011010110011101101011110100000" when "0111110011",
      "0101111111001001010111101101011001110011" when "0111110100",
      "0101111111110111111111101101010101000110" when "0111110101",
      "0110000000100110100111101101010000011000" when "0111110110",
      "0110000001010101001011101101001011101010" when "0111110111",
      "0110000010000011101111101101000110111011" when "0111111000",
      "0110000010110010010011101101000010001100" when "0111111001",
      "0110000011100000110011101100111101011011" when "0111111010",
      "0110000100001111010111101100111000101011" when "0111111011",
      "0110000100111101110111101100110011111010" when "0111111100",
      "0110000101101100010011101100101111001000" when "0111111101",
      "0110000110011010110011101100101010010110" when "0111111110",
      "0110000111001001001111101100100101100011" when "0111111111",
      "0110000111110111101111101100100000101111" when "1000000000",
      "0110001000100110000111101100011011111011" when "1000000001",
      "0110001001010100100011101100010111000110" when "1000000010",
      "0110001010000010111111101100010010010001" when "1000000011",
      "0110001010110001010111101100001101011011" when "1000000100",
      "0110001011011111101111101100001000100101" when "1000000101",
      "0110001100001110000011101100000011101110" when "1000000110",
      "0110001100111100011011101011111110110111" when "1000000111",
      "0110001101101010101111101011111001111111" when "1000001000",
      "0110001110011001000011101011110101000110" when "1000001001",
      "0110001111000111010111101011110000001101" when "1000001010",
      "0110001111110101100111101011101011010011" when "1000001011",
      "0110010000100011111011101011100110011001" when "1000001100",
      "0110010001010010001011101011100001011110" when "1000001101",
      "0110010010000000010111101011011100100011" when "1000001110",
      "0110010010101110100111101011010111100111" when "1000001111",
      "0110010011011100110011101011010010101010" when "1000010000",
      "0110010100001010111111101011001101101101" when "1000010001",
      "0110010100111001001011101011001000101111" when "1000010010",
      "0110010101100111010111101011000011110001" when "1000010011",
      "0110010110010101011111101010111110110010" when "1000010100",
      "0110010111000011100111101010111001110011" when "1000010101",
      "0110010111110001101111101010110100110011" when "1000010110",
      "0110011000011111110111101010101111110010" when "1000010111",
      "0110011001001101111011101010101010110001" when "1000011000",
      "0110011001111011111111101010100101101111" when "1000011001",
      "0110011010101010000011101010100000101101" when "1000011010",
      "0110011011011000000111101010011011101010" when "1000011011",
      "0110011100000110000111101010010110100111" when "1000011100",
      "0110011100110100000111101010010001100011" when "1000011101",
      "0110011101100010000111101010001100011110" when "1000011110",
      "0110011110010000000011101010000111011001" when "1000011111",
      "0110011110111110000011101010000010010100" when "1000100000",
      "0110011111101011111111101001111101001110" when "1000100001",
      "0110100000011001111011101001111000000111" when "1000100010",
      "0110100001000111110011101001110011000000" when "1000100011",
      "0110100001110101101111101001101101111000" when "1000100100",
      "0110100010100011100111101001101000101111" when "1000100101",
      "0110100011010001011111101001100011100110" when "1000100110",
      "0110100011111111010011101001011110011101" when "1000100111",
      "0110100100101101001011101001011001010010" when "1000101000",
      "0110100101011010111111101001010100001000" when "1000101001",
      "0110100110001000110011101001001110111101" when "1000101010",
      "0110100110110110100011101001001001110001" when "1000101011",
      "0110100111100100010111101001000100100100" when "1000101100",
      "0110101000010010000111101000111111010111" when "1000101101",
      "0110101000111111110011101000111010001010" when "1000101110",
      "0110101001101101100011101000110100111100" when "1000101111",
      "0110101010011011001111101000101111101101" when "1000110000",
      "0110101011001000111011101000101010011110" when "1000110001",
      "0110101011110110100111101000100101001110" when "1000110010",
      "0110101100100100010011101000011111111110" when "1000110011",
      "0110101101010001111011101000011010101101" when "1000110100",
      "0110101101111111100011101000010101011100" when "1000110101",
      "0110101110101101001011101000010000001010" when "1000110110",
      "0110101111011010101111101000001010110111" when "1000110111",
      "0110110000001000010111101000000101100100" when "1000111000",
      "0110110000110101111011101000000000010000" when "1000111001",
      "0110110001100011011011100111111010111100" when "1000111010",
      "0110110010010000111111100111110101100111" when "1000111011",
      "0110110010111110011111100111110000010010" when "1000111100",
      "0110110011101011111111100111101010111100" when "1000111101",
      "0110110100011001011111100111100101100110" when "1000111110",
      "0110110101000110111011100111100000001111" when "1000111111",
      "0110110101110100010111100111011010110111" when "1001000000",
      "0110110110100001110011100111010101011111" when "1001000001",
      "0110110111001111001111100111010000000110" when "1001000010",
      "0110110111111100100111100111001010101101" when "1001000011",
      "0110111000101001111111100111000101010011" when "1001000100",
      "0110111001010111010111100110111111111001" when "1001000101",
      "0110111010000100101111100110111010011110" when "1001000110",
      "0110111010110010000011100110110101000010" when "1001000111",
      "0110111011011111010111100110101111100110" when "1001001000",
      "0110111100001100101011100110101010001010" when "1001001001",
      "0110111100111001111011100110100100101101" when "1001001010",
      "0110111101100111001011100110011111001111" when "1001001011",
      "0110111110010100011011100110011001110001" when "1001001100",
      "0110111111000001101011100110010100010010" when "1001001101",
      "0110111111101110110111100110001110110010" when "1001001110",
      "0111000000011100000111100110001001010011" when "1001001111",
      "0111000001001001001111100110000011110010" when "1001010000",
      "0111000001110110011011100101111110010001" when "1001010001",
      "0111000010100011100011100101111000101111" when "1001010010",
      "0111000011010000101011100101110011001101" when "1001010011",
      "0111000011111101110011100101101101101011" when "1001010100",
      "0111000100101010111011100101101000000111" when "1001010101",
      "0111000101010111111111100101100010100100" when "1001010110",
      "0111000110000101000011100101011100111111" when "1001010111",
      "0111000110110010000111100101010111011010" when "1001011000",
      "0111000111011111000111100101010001110101" when "1001011001",
      "0111001000001100000111100101001100001111" when "1001011010",
      "0111001000111001000111100101000110101000" when "1001011011",
      "0111001001100110000111100101000001000001" when "1001011100",
      "0111001010010011000011100100111011011010" when "1001011101",
      "0111001010111111111111100100110101110001" when "1001011110",
      "0111001011101100111011100100110000001001" when "1001011111",
      "0111001100011001110011100100101010011111" when "1001100000",
      "0111001101000110101111100100100100110101" when "1001100001",
      "0111001101110011100111100100011111001011" when "1001100010",
      "0111001110100000011011100100011001100000" when "1001100011",
      "0111001111001101010011100100010011110100" when "1001100100",
      "0111001111111010000111100100001110001000" when "1001100101",
      "0111010000100110111011100100001000011100" when "1001100110",
      "0111010001010011101011100100000010101111" when "1001100111",
      "0111010010000000011011100011111101000001" when "1001101000",
      "0111010010101101001011100011110111010011" when "1001101001",
      "0111010011011001111011100011110001100100" when "1001101010",
      "0111010100000110101011100011101011110100" when "1001101011",
      "0111010100110011010111100011100110000101" when "1001101100",
      "0111010101100000000011100011100000010100" when "1001101101",
      "0111010110001100101011100011011010100011" when "1001101110",
      "0111010110111001010011100011010100110010" when "1001101111",
      "0111010111100101111011100011001110111111" when "1001110000",
      "0111011000010010100011100011001001001101" when "1001110001",
      "0111011000111111001011100011000011011010" when "1001110010",
      "0111011001101011101111100010111101100110" when "1001110011",
      "0111011010011000010011100010110111110001" when "1001110100",
      "0111011011000100110011100010110001111101" when "1001110101",
      "0111011011110001010111100010101100000111" when "1001110110",
      "0111011100011101110111100010100110010001" when "1001110111",
      "0111011101001010010011100010100000011011" when "1001111000",
      "0111011101110110110011100010011010100100" when "1001111001",
      "0111011110100011001111100010010100101100" when "1001111010",
      "0111011111001111101011100010001110110100" when "1001111011",
      "0111011111111100000011100010001000111011" when "1001111100",
      "0111100000101000011111100010000011000010" when "1001111101",
      "0111100001010100110111100001111101001001" when "1001111110",
      "0111100010000001001011100001110111001110" when "1001111111",
      "0111100010101101100011100001110001010011" when "1010000000",
      "0111100011011001110111100001101011011000" when "1010000001",
      "0111100100000110001011100001100101011100" when "1010000010",
      "0111100100110010011011100001011111100000" when "1010000011",
      "0111100101011110101111100001011001100011" when "1010000100",
      "0111100110001010111011100001010011100101" when "1010000101",
      "0111100110110111001011100001001101100111" when "1010000110",
      "0111100111100011011011100001000111101000" when "1010000111",
      "0111101000001111100111100001000001101001" when "1010001000",
      "0111101000111011101111100000111011101001" when "1010001001",
      "0111101001100111111011100000110101101001" when "1010001010",
      "0111101010010100000011100000101111101000" when "1010001011",
      "0111101011000000001011100000101001100111" when "1010001100",
      "0111101011101100010011100000100011100101" when "1010001101",
      "0111101100011000010111100000011101100011" when "1010001110",
      "0111101101000100011011100000010111100000" when "1010001111",
      "0111101101110000011111100000010001011100" when "1010010000",
      "0111101110011100011111100000001011011000" when "1010010001",
      "0111101111001000011111100000000101010011" when "1010010010",
      "0111101111110100011111011111111111001110" when "1010010011",
      "0111110000100000011011011111111001001001" when "1010010100",
      "0111110001001100011011011111110011000010" when "1010010101",
      "0111110001111000010111011111101100111100" when "1010010110",
      "0111110010100100001111011111100110110100" when "1010010111",
      "0111110011010000001011011111100000101100" when "1010011000",
      "0111110011111100000011011111011010100100" when "1010011001",
      "0111110100100111110111011111010100011011" when "1010011010",
      "0111110101010011101111011111001110010010" when "1010011011",
      "0111110101111111100011011111001000001000" when "1010011100",
      "0111110110101011010111011111000001111101" when "1010011101",
      "0111110111010111000111011110111011110010" when "1010011110",
      "0111111000000010110111011110110101100111" when "1010011111",
      "0111111000101110100111011110101111011010" when "1010100000",
      "0111111001011010010111011110101001001110" when "1010100001",
      "0111111010000110000011011110100011000001" when "1010100010",
      "0111111010110001101111011110011100110011" when "1010100011",
      "0111111011011101011011011110010110100100" when "1010100100",
      "0111111100001001000011011110010000010110" when "1010100101",
      "0111111100110100101011011110001010000110" when "1010100110",
      "0111111101100000010011011110000011110110" when "1010100111",
      "0111111110001011111011011101111101100110" when "1010101000",
      "0111111110110111011111011101110111010101" when "1010101001",
      "0111111111100011000011011101110001000100" when "1010101010",
      "1000000000001110100011011101101010110010" when "1010101011",
      "1000000000111010000011011101100100011111" when "1010101100",
      "1000000001100101100011011101011110001100" when "1010101101",
      "1000000010010001000011011101010111111000" when "1010101110",
      "1000000010111100011111011101010001100100" when "1010101111",
      "1000000011100111111011011101001011001111" when "1010110000",
      "1000000100010011010111011101000100111010" when "1010110001",
      "1000000100111110101111011100111110100100" when "1010110010",
      "1000000101101010000111011100111000001110" when "1010110011",
      "1000000110010101011111011100110001110111" when "1010110100",
      "1000000111000000110111011100101011100000" when "1010110101",
      "1000000111101100001011011100100101001000" when "1010110110",
      "1000001000010111011011011100011110110000" when "1010110111",
      "1000001001000010101111011100011000010111" when "1010111000",
      "1000001001101101111111011100010001111101" when "1010111001",
      "1000001010011001001111011100001011100011" when "1010111010",
      "1000001011000100011111011100000101001001" when "1010111011",
      "1000001011101111101011011011111110101110" when "1010111100",
      "1000001100011010110111011011111000010010" when "1010111101",
      "1000001101000101111111011011110001110110" when "1010111110",
      "1000001101110001001011011011101011011001" when "1010111111",
      "1000001110011100010011011011100100111100" when "1011000000",
      "1000001111000111010111011011011110011110" when "1011000001",
      "1000001111110010011111011011011000000000" when "1011000010",
      "1000010000011101100011011011010001100001" when "1011000011",
      "1000010001001000100011011011001011000010" when "1011000100",
      "1000010001110011100111011011000100100010" when "1011000101",
      "1000010010011110100111011010111110000010" when "1011000110",
      "1000010011001001100011011010110111100001" when "1011000111",
      "1000010011110100100011011010110000111111" when "1011001000",
      "1000010100011111011111011010101010011101" when "1011001001",
      "1000010101001010011011011010100011111011" when "1011001010",
      "1000010101110101010011011010011101011000" when "1011001011",
      "1000010110100000001011011010010110110100" when "1011001100",
      "1000010111001011000011011010010000010000" when "1011001101",
      "1000010111110101111011011010001001101100" when "1011001110",
      "1000011000100000101111011010000011000111" when "1011001111",
      "1000011001001011100011011001111100100001" when "1011010000",
      "1000011001110110010011011001110101111011" when "1011010001",
      "1000011010100001000011011001101111010100" when "1011010010",
      "1000011011001011110011011001101000101101" when "1011010011",
      "1000011011110110100011011001100010000101" when "1011010100",
      "1000011100100001001111011001011011011101" when "1011010101",
      "1000011101001011111011011001010100110100" when "1011010110",
      "1000011101110110100111011001001110001011" when "1011010111",
      "1000011110100001001111011001000111100001" when "1011011000",
      "1000011111001011110111011001000000110111" when "1011011001",
      "1000011111110110011011011000111010001100" when "1011011010",
      "1000100000100001000011011000110011100000" when "1011011011",
      "1000100001001011100111011000101100110101" when "1011011100",
      "1000100001110110000111011000100110001000" when "1011011101",
      "1000100010100000101011011000011111011011" when "1011011110",
      "1000100011001011000111011000011000101110" when "1011011111",
      "1000100011110101100111011000010010000000" when "1011100000",
      "1000100100100000000011011000001011010001" when "1011100001",
      "1000100101001010011111011000000100100010" when "1011100010",
      "1000100101110100111011010111111101110011" when "1011100011",
      "1000100110011111010011010111110111000010" when "1011100100",
      "1000100111001001101011010111110000010010" when "1011100101",
      "1000100111110100000011010111101001100001" when "1011100110",
      "1000101000011110010111010111100010101111" when "1011100111",
      "1000101001001000101011010111011011111101" when "1011101000",
      "1000101001110010111111010111010101001010" when "1011101001",
      "1000101010011101001111010111001110010111" when "1011101010",
      "1000101011000111011111010111000111100011" when "1011101011",
      "1000101011110001101111010111000000101111" when "1011101100",
      "1000101100011011111011010110111001111010" when "1011101101",
      "1000101101000110000111010110110011000101" when "1011101110",
      "1000101101110000010011010110101100001111" when "1011101111",
      "1000101110011010011011010110100101011001" when "1011110000",
      "1000101111000100100011010110011110100010" when "1011110001",
      "1000101111101110101011010110010111101011" when "1011110010",
      "1000110000011000101111010110010000110011" when "1011110011",
      "1000110001000010110011010110001001111010" when "1011110100",
      "1000110001101100110011010110000011000010" when "1011110101",
      "1000110010010110110111010101111100001000" when "1011110110",
      "1000110011000000110111010101110101001110" when "1011110111",
      "1000110011101010110011010101101110010100" when "1011111000",
      "1000110100010100101111010101100111011001" when "1011111001",
      "1000110100111110101011010101100000011101" when "1011111010",
      "1000110101101000100111010101011001100001" when "1011111011",
      "1000110110010010011111010101010010100101" when "1011111100",
      "1000110110111100010111010101001011101000" when "1011111101",
      "1000110111100110001111010101000100101010" when "1011111110",
      "1000111000010000000011010100111101101100" when "1011111111",
      "1000111000111001110111010100110110101110" when "1100000000",
      "1000111001100011100111010100101111101111" when "1100000001",
      "1000111010001101010111010100101000101111" when "1100000010",
      "1000111010110111000111010100100001101111" when "1100000011",
      "1000111011100000110111010100011010101110" when "1100000100",
      "1000111100001010100011010100010011101101" when "1100000101",
      "1000111100110100001111010100001100101100" when "1100000110",
      "1000111101011101110111010100000101101010" when "1100000111",
      "1000111110000111011111010011111110100111" when "1100001000",
      "1000111110110001000111010011110111100100" when "1100001001",
      "1000111111011010101011010011110000100000" when "1100001010",
      "1001000000000100010011010011101001011100" when "1100001011",
      "1001000000101101110011010011100010010111" when "1100001100",
      "1001000001010111010111010011011011010010" when "1100001101",
      "1001000010000000110111010011010100001100" when "1100001110",
      "1001000010101010010011010011001101000110" when "1100001111",
      "1001000011010011110011010011000101111111" when "1100010000",
      "1001000011111101001111010010111110111000" when "1100010001",
      "1001000100100110100111010010110111110000" when "1100010010",
      "1001000101010000000011010010110000101000" when "1100010011",
      "1001000101111001011011010010101001011111" when "1100010100",
      "1001000110100010101111010010100010010110" when "1100010101",
      "1001000111001100000011010010011011001100" when "1100010110",
      "1001000111110101010111010010010100000010" when "1100010111",
      "1001001000011110101011010010001100110111" when "1100011000",
      "1001001001000111111011010010000101101100" when "1100011001",
      "1001001001110001001011010001111110100000" when "1100011010",
      "1001001010011010010111010001110111010100" when "1100011011",
      "1001001011000011100011010001110000000111" when "1100011100",
      "1001001011101100101111010001101000111010" when "1100011101",
      "1001001100010101111011010001100001101100" when "1100011110",
      "1001001100111111000011010001011010011110" when "1100011111",
      "1001001101101000000111010001010011001111" when "1100100000",
      "1001001110010001001111010001001011111111" when "1100100001",
      "1001001110111010010011010001000100110000" when "1100100010",
      "1001001111100011010011010000111101011111" when "1100100011",
      "1001010000001100010111010000110110001110" when "1100100100",
      "1001010000110101010111010000101110111101" when "1100100101",
      "1001010001011110010011010000100111101011" when "1100100110",
      "1001010010000111001111010000100000011001" when "1100100111",
      "1001010010110000001011010000011001000110" when "1100101000",
      "1001010011011001000111010000010001110011" when "1100101001",
      "1001010100000001111111010000001010011111" when "1100101010",
      "1001010100101010110111010000000011001010" when "1100101011",
      "1001010101010011101011001111111011110101" when "1100101100",
      "1001010101111100011111001111110100100000" when "1100101101",
      "1001010110100101010011001111101101001010" when "1100101110",
      "1001010111001110000011001111100101110100" when "1100101111",
      "1001010111110110110011001111011110011101" when "1100110000",
      "1001011000011111100011001111010111000110" when "1100110001",
      "1001011001001000001111001111001111101110" when "1100110010",
      "1001011001110000111011001111001000010101" when "1100110011",
      "1001011010011001100111001111000000111101" when "1100110100",
      "1001011011000010001111001110111001100011" when "1100110101",
      "1001011011101010110011001110110010001001" when "1100110110",
      "1001011100010011011011001110101010101111" when "1100110111",
      "1001011100111011111111001110100011010100" when "1100111000",
      "1001011101100100100011001110011011111001" when "1100111001",
      "1001011110001101000011001110010100011101" when "1100111010",
      "1001011110110101100011001110001101000001" when "1100111011",
      "1001011111011110000011001110000101100100" when "1100111100",
      "1001100000000110011111001101111110000110" when "1100111101",
      "1001100000101110111011001101110110101000" when "1100111110",
      "1001100001010111010011001101101111001010" when "1100111111",
      "1001100001111111101011001101100111101011" when "1101000000",
      "1001100010101000000011001101100000001100" when "1101000001",
      "1001100011010000011011001101011000101100" when "1101000010",
      "1001100011111000101111001101010001001100" when "1101000011",
      "1001100100100000111111001101001001101011" when "1101000100",
      "1001100101001001010011001101000010001010" when "1101000101",
      "1001100101110001100011001100111010101000" when "1101000110",
      "1001100110011001101111001100110011000110" when "1101000111",
      "1001100111000001111011001100101011100011" when "1101001000",
      "1001100111101010000111001100100100000000" when "1101001001",
      "1001101000010010010011001100011100011100" when "1101001010",
      "1001101000111010011011001100010100110111" when "1101001011",
      "1001101001100010100011001100001101010011" when "1101001100",
      "1001101010001010100111001100000101101101" when "1101001101",
      "1001101010110010101011001011111110001000" when "1101001110",
      "1001101011011010101011001011110110100001" when "1101001111",
      "1001101100000010101111001011101110111011" when "1101010000",
      "1001101100101010101111001011100111010100" when "1101010001",
      "1001101101010010101011001011011111101100" when "1101010010",
      "1001101101111010100111001011011000000100" when "1101010011",
      "1001101110100010100011001011010000011011" when "1101010100",
      "1001101111001010011011001011001000110010" when "1101010101",
      "1001101111110010010011001011000001001000" when "1101010110",
      "1001110000011010001011001010111001011110" when "1101010111",
      "1001110001000001111111001010110001110011" when "1101011000",
      "1001110001101001110011001010101010001000" when "1101011001",
      "1001110010010001100011001010100010011101" when "1101011010",
      "1001110010111001010011001010011010110000" when "1101011011",
      "1001110011100001000011001010010011000100" when "1101011100",
      "1001110100001000101111001010001011010111" when "1101011101",
      "1001110100110000011011001010000011101001" when "1101011110",
      "1001110101011000000111001001111011111011" when "1101011111",
      "1001110101111111101111001001110100001101" when "1101100000",
      "1001110110100111010111001001101100011101" when "1101100001",
      "1001110111001110111111001001100100101110" when "1101100010",
      "1001110111110110100011001001011100111110" when "1101100011",
      "1001111000011110000011001001010101001101" when "1101100100",
      "1001111001000101100111001001001101011101" when "1101100101",
      "1001111001101101000011001001000101101011" when "1101100110",
      "1001111010010100100011001000111101111001" when "1101100111",
      "1001111010111011111111001000110110000111" when "1101101000",
      "1001111011100011011011001000101110010100" when "1101101001",
      "1001111100001010110011001000100110100000" when "1101101010",
      "1001111100110010001011001000011110101100" when "1101101011",
      "1001111101011001100011001000010110111000" when "1101101100",
      "1001111110000000110111001000001111000011" when "1101101101",
      "1001111110101000001011001000000111001110" when "1101101110",
      "1001111111001111011111000111111111011000" when "1101101111",
      "1001111111110110101111000111110111100010" when "1101110000",
      "1010000000011101111011000111101111101011" when "1101110001",
      "1010000001000101001011000111100111110100" when "1101110010",
      "1010000001101100010111000111011111111100" when "1101110011",
      "1010000010010011011111000111011000000100" when "1101110100",
      "1010000010111010100111000111010000001011" when "1101110101",
      "1010000011100001101111000111001000010010" when "1101110110",
      "1010000100001000110011000111000000011000" when "1101110111",
      "1010000100101111110111000110111000011110" when "1101111000",
      "1010000101010110111011000110110000100100" when "1101111001",
      "1010000101111101111011000110101000101000" when "1101111010",
      "1010000110100100111011000110100000101101" when "1101111011",
      "1010000111001011111011000110011000110001" when "1101111100",
      "1010000111110010110111000110010000110100" when "1101111101",
      "1010001000011001101111000110001000110111" when "1101111110",
      "1010001001000000101011000110000000111010" when "1101111111",
      "1010001001100111011111000101111000111100" when "1110000000",
      "1010001010001110010111000101110000111101" when "1110000001",
      "1010001010110101001011000101101000111110" when "1110000010",
      "1010001011011011111111000101100000111111" when "1110000011",
      "1010001100000010101111000101011000111111" when "1110000100",
      "1010001100101001011111000101010000111111" when "1110000101",
      "1010001101010000001011000101001000111110" when "1110000110",
      "1010001101110110111011000101000000111101" when "1110000111",
      "1010001110011101100011000100111000111011" when "1110001000",
      "1010001111000100001111000100110000111001" when "1110001001",
      "1010001111101010110111000100101000110110" when "1110001010",
      "1010010000010001011011000100100000110011" when "1110001011",
      "1010010000110111111111000100011000101111" when "1110001100",
      "1010010001011110100011000100010000101011" when "1110001101",
      "1010010010000101000011000100001000100110" when "1110001110",
      "1010010010101011100011000100000000100001" when "1110001111",
      "1010010011010010000011000011111000011100" when "1110010000",
      "1010010011111000011111000011110000010110" when "1110010001",
      "1010010100011110111011000011101000001111" when "1110010010",
      "1010010101000101010011000011100000001000" when "1110010011",
      "1010010101101011101011000011011000000001" when "1110010100",
      "1010010110010010000011000011001111111001" when "1110010101",
      "1010010110111000010111000011000111110001" when "1110010110",
      "1010010111011110101011000010111111101000" when "1110010111",
      "1010011000000100111011000010110111011110" when "1110011000",
      "1010011000101011001011000010101111010101" when "1110011001",
      "1010011001010001011011000010100111001010" when "1110011010",
      "1010011001110111100111000010011111000000" when "1110011011",
      "1010011010011101110011000010010110110100" when "1110011100",
      "1010011011000011111011000010001110101001" when "1110011101",
      "1010011011101010000011000010000110011101" when "1110011110",
      "1010011100010000001011000001111110010000" when "1110011111",
      "1010011100110110001111000001110110000011" when "1110100000",
      "1010011101011100010011000001101101110101" when "1110100001",
      "1010011110000010010011000001100101100111" when "1110100010",
      "1010011110101000010011000001011101011001" when "1110100011",
      "1010011111001110010011000001010101001010" when "1110100100",
      "1010011111110100001111000001001100111011" when "1110100101",
      "1010100000011010000111000001000100101011" when "1110100110",
      "1010100001000000000011000000111100011010" when "1110100111",
      "1010100001100101111011000000110100001010" when "1110101000",
      "1010100010001011101111000000101011111000" when "1110101001",
      "1010100010110001100011000000100011100111" when "1110101010",
      "1010100011010111010111000000011011010100" when "1110101011",
      "1010100011111101000111000000010011000010" when "1110101100",
      "1010100100100010110111000000001010101111" when "1110101101",
      "1010100101001000100111000000000010011011" when "1110101110",
      "1010100101101110010010111111111010000111" when "1110101111",
      "1010100110010011111110111111110001110010" when "1110110000",
      "1010100110111001100110111111101001011101" when "1110110001",
      "1010100111011111001110111111100001001000" when "1110110010",
      "1010101000000100110010111111011000110010" when "1110110011",
      "1010101000101010010110111111010000011100" when "1110110100",
      "1010101001001111111010111111001000000101" when "1110110101",
      "1010101001110101011010111110111111101110" when "1110110110",
      "1010101010011010111010111110110111010110" when "1110110111",
      "1010101011000000010110111110101110111110" when "1110111000",
      "1010101011100101110010111110100110100101" when "1110111001",
      "1010101100001011001110111110011110001100" when "1110111010",
      "1010101100110000100110111110010101110010" when "1110111011",
      "1010101101010101111110111110001101011000" when "1110111100",
      "1010101101111011010010111110000100111110" when "1110111101",
      "1010101110100000100110111101111100100011" when "1110111110",
      "1010101111000101111010111101110100001000" when "1110111111",
      "1010101111101011001010111101101011101100" when "1111000000",
      "1010110000010000011010111101100011001111" when "1111000001",
      "1010110000110101100110111101011010110011" when "1111000010",
      "1010110001011010110010111101010010010101" when "1111000011",
      "1010110001111111111010111101001001111000" when "1111000100",
      "1010110010100101000010111101000001011010" when "1111000101",
      "1010110011001010001010111100111000111011" when "1111000110",
      "1010110011101111001110111100110000011100" when "1111000111",
      "1010110100010100010010111100100111111100" when "1111001000",
      "1010110100111001010010111100011111011100" when "1111001001",
      "1010110101011110010010111100010110111100" when "1111001010",
      "1010110110000011010010111100001110011011" when "1111001011",
      "1010110110101000001110111100000101111010" when "1111001100",
      "1010110111001101000110111011111101011000" when "1111001101",
      "1010110111110010000010111011110100110110" when "1111001110",
      "1010111000010110111010111011101100010011" when "1111001111",
      "1010111000111011101110111011100011110000" when "1111010000",
      "1010111001100000100010111011011011001100" when "1111010001",
      "1010111010000101010110111011010010101000" when "1111010010",
      "1010111010101010000110111011001010000100" when "1111010011",
      "1010111011001110110110111011000001011111" when "1111010100",
      "1010111011110011100010111010111000111010" when "1111010101",
      "1010111100011000001110111010110000010100" when "1111010110",
      "1010111100111100110110111010100111101101" when "1111010111",
      "1010111101100001011110111010011111000111" when "1111011000",
      "1010111110000110000110111010010110011111" when "1111011001",
      "1010111110101010101010111010001101111000" when "1111011010",
      "1010111111001111001110111010000101010000" when "1111011011",
      "1010111111110011101110111001111100100111" when "1111011100",
      "1011000000011000001110111001110011111110" when "1111011101",
      "1011000000111100101110111001101011010101" when "1111011110",
      "1011000001100001001010111001100010101011" when "1111011111",
      "1011000010000101100110111001011010000001" when "1111100000",
      "1011000010101001111110111001010001010110" when "1111100001",
      "1011000011001110010110111001001000101011" when "1111100010",
      "1011000011110010101010111000111111111111" when "1111100011",
      "1011000100010110111110111000110111010011" when "1111100100",
      "1011000100111011010010111000101110100110" when "1111100101",
      "1011000101011111100010111000100101111001" when "1111100110",
      "1011000110000011101110111000011101001100" when "1111100111",
      "1011000110100111111110111000010100011110" when "1111101000",
      "1011000111001100001010111000001011101111" when "1111101001",
      "1011000111110000010010111000000011000001" when "1111101010",
      "1011001000010100011010110111111010010001" when "1111101011",
      "1011001000111000011110110111110001100010" when "1111101100",
      "1011001001011100100110110111101000110010" when "1111101101",
      "1011001010000000100110110111100000000001" when "1111101110",
      "1011001010100100101010110111010111010000" when "1111101111",
      "1011001011001000100110110111001110011111" when "1111110000",
      "1011001011101100100110110111000101101101" when "1111110001",
      "1011001100010000100010110110111100111011" when "1111110010",
      "1011001100110100011010110110110100001000" when "1111110011",
      "1011001101011000010010110110101011010101" when "1111110100",
      "1011001101111100001010110110100010100001" when "1111110101",
      "1011001110011111111110110110011001101101" when "1111110110",
      "1011001111000011110010110110010000111000" when "1111110111",
      "1011001111100111100110110110001000000011" when "1111111000",
      "1011010000001011010010110101111111001110" when "1111111001",
      "1011010000101111000010110101110110011000" when "1111111010",
      "1011010001010010101110110101101101100010" when "1111111011",
      "1011010001110110011010110101100100101011" when "1111111100",
      "1011010010011010000010110101011011110100" when "1111111101",
      "1011010010111101101010110101010010111100" when "1111111110",
      "1011010011100001001110110101001010000100" when "1111111111",
      "----------------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_10_comb_uid14
-- VHDL generated for Virtex6 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: 1.021000nsY: 1.021000nsCin: 0.000000ns
--  approx. output signal timings: R: 1.921000ns

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_10_comb_uid14 is
    port (X : in  std_logic_vector(9 downto 0);
          Y : in  std_logic_vector(9 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(9 downto 0)   );
end entity;

architecture arch of IntAdder_10_comb_uid14 is
signal Rtmp :  std_logic_vector(9 downto 0);
   -- timing of Rtmp: 1.921000ns
begin
   Rtmp <= X + Y + Cin;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                            FixRealKCM_comb_uid6
-- VHDL generated for Virtex6 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: 0.366000ns
--  approx. output signal timings: R: 1.921000ns

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_comb_uid6 is
    port (X : in  std_logic_vector(7 downto 0);
          R : out  std_logic_vector(9 downto 0)   );
end entity;

architecture arch of FixRealKCM_comb_uid6 is
   component FixRealKCM_comb_uid6_T0_comb_uid9 is
      port ( X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(9 downto 0)   );
   end component;

   component FixRealKCM_comb_uid6_T1_comb_uid11 is
      port ( X : in  std_logic_vector(1 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntAdder_10_comb_uid14 is
      port ( X : in  std_logic_vector(9 downto 0);
             Y : in  std_logic_vector(9 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(9 downto 0)   );
   end component;

signal FixRealKCM_comb_uid6_A0 :  std_logic_vector(5 downto 0);
   -- timing of FixRealKCM_comb_uid6_A0: 0.366000ns
signal FixRealKCM_comb_uid6_T0 :  std_logic_vector(9 downto 0);
   -- timing of FixRealKCM_comb_uid6_T0: 1.021000ns
signal bh7_w0_0 :  std_logic;
   -- timing of bh7_w0_0: 1.021000ns
signal bh7_w1_0 :  std_logic;
   -- timing of bh7_w1_0: 1.021000ns
signal bh7_w2_0 :  std_logic;
   -- timing of bh7_w2_0: 1.021000ns
signal bh7_w3_0 :  std_logic;
   -- timing of bh7_w3_0: 1.021000ns
signal bh7_w4_0 :  std_logic;
   -- timing of bh7_w4_0: 1.021000ns
signal bh7_w5_0 :  std_logic;
   -- timing of bh7_w5_0: 1.021000ns
signal bh7_w6_0 :  std_logic;
   -- timing of bh7_w6_0: 1.021000ns
signal bh7_w7_0 :  std_logic;
   -- timing of bh7_w7_0: 1.021000ns
signal bh7_w8_0 :  std_logic;
   -- timing of bh7_w8_0: 1.021000ns
signal bh7_w9_0 :  std_logic;
   -- timing of bh7_w9_0: 1.021000ns
signal FixRealKCM_comb_uid6_A1 :  std_logic_vector(1 downto 0);
   -- timing of FixRealKCM_comb_uid6_A1: 0.366000ns
signal FixRealKCM_comb_uid6_T1 :  std_logic_vector(3 downto 0);
   -- timing of FixRealKCM_comb_uid6_T1: 1.015000ns
signal bh7_w0_1 :  std_logic;
   -- timing of bh7_w0_1: 1.015000ns
signal bh7_w1_1 :  std_logic;
   -- timing of bh7_w1_1: 1.015000ns
signal bh7_w2_1 :  std_logic;
   -- timing of bh7_w2_1: 1.015000ns
signal bh7_w3_1 :  std_logic;
   -- timing of bh7_w3_1: 1.015000ns
signal bitheapFinalAdd_bh7_In0 :  std_logic_vector(9 downto 0);
   -- timing of bitheapFinalAdd_bh7_In0: 1.021000ns
signal bitheapFinalAdd_bh7_In1 :  std_logic_vector(9 downto 0);
   -- timing of bitheapFinalAdd_bh7_In1: 1.021000ns
signal bitheapFinalAdd_bh7_Cin :  std_logic;
   -- timing of bitheapFinalAdd_bh7_Cin: 0.000000ns
signal bitheapFinalAdd_bh7_Out :  std_logic_vector(9 downto 0);
   -- timing of bitheapFinalAdd_bh7_Out: 1.921000ns
signal bitheapResult_bh7 :  std_logic_vector(9 downto 0);
   -- timing of bitheapResult_bh7: 1.921000ns
signal OutRes :  std_logic_vector(9 downto 0);
   -- timing of OutRes: 1.921000ns
begin
-- This operator multiplies by pi
   FixRealKCM_comb_uid6_A0 <= X(7 downto 2);-- input address  m=-13  l=-18
   FixRealKCM_comb_uid6_Table0: FixRealKCM_comb_uid6_T0_comb_uid9
      port map ( X => FixRealKCM_comb_uid6_A0,
                 Y => FixRealKCM_comb_uid6_T0);
   bh7_w0_0 <= FixRealKCM_comb_uid6_T0(0);
   bh7_w1_0 <= FixRealKCM_comb_uid6_T0(1);
   bh7_w2_0 <= FixRealKCM_comb_uid6_T0(2);
   bh7_w3_0 <= FixRealKCM_comb_uid6_T0(3);
   bh7_w4_0 <= FixRealKCM_comb_uid6_T0(4);
   bh7_w5_0 <= FixRealKCM_comb_uid6_T0(5);
   bh7_w6_0 <= FixRealKCM_comb_uid6_T0(6);
   bh7_w7_0 <= FixRealKCM_comb_uid6_T0(7);
   bh7_w8_0 <= FixRealKCM_comb_uid6_T0(8);
   bh7_w9_0 <= FixRealKCM_comb_uid6_T0(9);
   FixRealKCM_comb_uid6_A1 <= X(1 downto 0);-- input address  m=-19  l=-20
   FixRealKCM_comb_uid6_Table1: FixRealKCM_comb_uid6_T1_comb_uid11
      port map ( X => FixRealKCM_comb_uid6_A1,
                 Y => FixRealKCM_comb_uid6_T1);
   bh7_w0_1 <= FixRealKCM_comb_uid6_T1(0);
   bh7_w1_1 <= FixRealKCM_comb_uid6_T1(1);
   bh7_w2_1 <= FixRealKCM_comb_uid6_T1(2);
   bh7_w3_1 <= FixRealKCM_comb_uid6_T1(3);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   bitheapFinalAdd_bh7_In0 <= "" & bh7_w9_0 & bh7_w8_0 & bh7_w7_0 & bh7_w6_0 & bh7_w5_0 & bh7_w4_0 & bh7_w3_1 & bh7_w2_1 & bh7_w1_1 & bh7_w0_1;
   bitheapFinalAdd_bh7_In1 <= "0" & "0" & "0" & "0" & "0" & "0" & bh7_w3_0 & bh7_w2_0 & bh7_w1_0 & bh7_w0_0;
   bitheapFinalAdd_bh7_Cin <= '0';

   bitheapFinalAdd_bh7: IntAdder_10_comb_uid14
      port map ( Cin => bitheapFinalAdd_bh7_Cin,
                 X => bitheapFinalAdd_bh7_In0,
                 Y => bitheapFinalAdd_bh7_In1,
                 R => bitheapFinalAdd_bh7_Out);
   bitheapResult_bh7 <= bitheapFinalAdd_bh7_Out(9 downto 0);
   OutRes <= bitheapResult_bh7(9 downto 0);
   R <= OutRes(9 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                       FixSinCosPoly_LSBm16_comb_uid2
-- VHDL generated for Virtex6 @ 0MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Antoine Martinet, Guillaume Sergent, (2013-2019)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): inf
-- Target frequency (MHz): 0
-- Input signals: X
-- Output signals: S C
--  approx. input signal timings: X: 0.000000ns
--  approx. output signal timings: S: 4.924000nsC: 4.924000ns

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixSinCosPoly_LSBm16_comb_uid2 is
    port (X : in  std_logic_vector(16 downto 0);
          S : out  std_logic_vector(16 downto 0);
          C : out  std_logic_vector(16 downto 0)   );
end entity;

architecture arch of FixSinCosPoly_LSBm16_comb_uid2 is
   component SinCosTable_comb_uid4 is
      port ( X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(39 downto 0)   );
   end component;

   component FixRealKCM_comb_uid6 is
      port ( X : in  std_logic_vector(7 downto 0);
             R : out  std_logic_vector(9 downto 0)   );
   end component;

signal X_sgn :  std_logic;
   -- timing of X_sgn: 0.000000ns
signal Q :  std_logic;
   -- timing of Q: 0.000000ns
signal O :  std_logic;
   -- timing of O: 0.000000ns
signal Y :  std_logic_vector(13 downto 0);
   -- timing of Y: 0.000000ns
signal Yneg :  std_logic_vector(17 downto 0);
   -- timing of Yneg: 0.366000ns
signal A :  std_logic_vector(9 downto 0);
   -- timing of A: 0.366000ns
signal Y_red :  std_logic_vector(7 downto 0);
   -- timing of Y_red: 0.366000ns
signal SinCosA :  std_logic_vector(39 downto 0);
   -- timing of SinCosA: 2.236000ns
signal SinPiA :  std_logic_vector(19 downto 0);
   -- timing of SinPiA: 2.236000ns
signal CosPiA :  std_logic_vector(19 downto 0);
   -- timing of CosPiA: 2.236000ns
signal Z :  std_logic_vector(9 downto 0);
   -- timing of Z: 1.921000ns
signal SinPiACosZ :  std_logic_vector(19 downto 0);
   -- timing of SinPiACosZ: 2.236000ns
signal CosPiAtrunc :  std_logic_vector(9 downto 0);
   -- timing of CosPiAtrunc: 2.236000ns
signal CosPiASinZ :  std_logic_vector(19 downto 0);
   -- timing of CosPiASinZ: 3.874000ns
signal PreSinX :  std_logic_vector(19 downto 0);
   -- timing of PreSinX: 4.924000ns
signal CosPiACosZ :  std_logic_vector(19 downto 0);
   -- timing of CosPiACosZ: 2.236000ns
signal SinPiAtrunc :  std_logic_vector(9 downto 0);
   -- timing of SinPiAtrunc: 2.236000ns
signal SinPiASinZ :  std_logic_vector(19 downto 0);
   -- timing of SinPiASinZ: 2.236000ns
signal PreCosX :  std_logic_vector(19 downto 0);
   -- timing of PreCosX: 3.286000ns
signal C_out :  std_logic_vector(15 downto 0);
   -- timing of C_out: 3.286000ns
signal S_out :  std_logic_vector(15 downto 0);
   -- timing of S_out: 4.924000ns
signal C_sgn :  std_logic;
   -- timing of C_sgn: 0.000000ns
signal Exch :  std_logic;
   -- timing of Exch: 0.000000ns
signal S_wo_sgn :  std_logic_vector(15 downto 0);
   -- timing of S_wo_sgn: 4.924000ns
signal C_wo_sgn :  std_logic_vector(15 downto 0);
   -- timing of C_wo_sgn: 4.924000ns
signal S_wo_sgn_ext :  std_logic_vector(16 downto 0);
   -- timing of S_wo_sgn_ext: 4.924000ns
signal C_wo_sgn_ext :  std_logic_vector(16 downto 0);
   -- timing of C_wo_sgn_ext: 4.924000ns
signal S_wo_sgn_neg :  std_logic_vector(16 downto 0);
   -- timing of S_wo_sgn_neg: 4.924000ns
signal C_wo_sgn_neg :  std_logic_vector(16 downto 0);
   -- timing of C_wo_sgn_neg: 4.924000ns
begin
   -- The argument is reduced into (0,1/4)
   X_sgn <= X(16);  -- sign
   Q <= X(15);  -- quadrant
   O <= X(14);  -- octant
   Y <= X (13 downto 0);
   -- Computing .25-Y :  we do a logic NOT, at a cost of 1 ulp
   Yneg <= ((not Y) & "1111") when O='1' else (Y & "0000");
   A <= Yneg (17 downto 8);
   Y_red <= Yneg(7 downto 0);
   SinCosTable: SinCosTable_comb_uid4
      port map ( X => A,
                 Y => SinCosA);
   SinPiA <= SinCosA(39 downto 20);
   CosPiA <= SinCosA(19 downto 0);
   MultByPi: FixRealKCM_comb_uid6
      port map ( X => Y_red,
                 R => Z);
   SinPiACosZ <= SinPiA; -- For these sizes  CosZ approx 1
   CosPiAtrunc <= CosPiA(19 downto 10);
   CosPiASinZ <= CosPiAtrunc*Z;  -- For these sizes  SinZ approx Z
   PreSinX <= SinPiACosZ + ( "0000000000" & (CosPiASinZ(19 downto 10)) );
   CosPiACosZ <= CosPiA; -- For these sizes  CosZ approx 1
   SinPiAtrunc <= SinPiA(19 downto 10);
   SinPiASinZ <= SinPiAtrunc*Z;  -- For these sizes  SinZ approx Z
   PreCosX <= CosPiACosZ - ( "0000000000" & (SinPiASinZ(19 downto 10)) );
   C_out <= PreCosX(19 downto 4);
   S_out <= PreSinX(19 downto 4);
   -- --- Final reconstruction of both sine and cosine ---
   C_sgn <= X_sgn xor Q;
   Exch <= Q xor O;
   S_wo_sgn <= C_out when Exch = '1' else S_out;
   C_wo_sgn <= S_out when Exch = '1' else C_out;
   S_wo_sgn_ext <= '0' & S_wo_sgn;
   C_wo_sgn_ext <= '0' & C_wo_sgn;
   S_wo_sgn_neg <= (not S_wo_sgn_ext) + 1;
   C_wo_sgn_neg <= (not C_wo_sgn_ext) + 1;
   S <= S_wo_sgn_ext when X_sgn = '0' else S_wo_sgn_neg;
   C <= C_wo_sgn_ext when C_sgn = '0' else C_wo_sgn_neg;
end architecture;

